
module johnson_counter(Clock,
    Reset,
    Count_out
    );
    input Clock;
    input Reset;
    output [3:0] Count_out;
    reg [3:0] Count_temp;
    always @(posedge(Clock) or Reset)
    begin
        if(Reset == 1'b1)   begin
            Count_temp = 4'b0000;   end
        else if(Clock == 1'b1)  begin
            Count_temp = {Count_temp[2:0],~Count_temp[3]};  end 
    end
    assign Count_out = Count_temp;
endmodule

module johnson_ring;
    reg Clock;
    reg Reset;
    wire [3:0] Count_out;
    johnson_counter uut (
        .Clock(Clock), 
        .Reset(Reset), 
        .Count_out(Count_out)
    );
    initial Clock = 0; 
    always #10 Clock = ~Clock;     
    initial begin
        Reset = 1; 
        #50;
        Reset = 0;
    end
      
endmodule